CONFIGURATION cfg OF contatore_tb IS
   FOR contatore_test
      -- use default configuration
   END FOR;
END cfg;
